module multiplier(
    input [15:0] a,
    input [15:0] b,
    output [31:0] answer
);


endmodule