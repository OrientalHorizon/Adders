module Booth(
    input   [15:0]  a,
    input   [15:0]  b,
    input           clk,
    output  [31:0]  mul
);

    wire [15:0] a_neg;
    assign a_neg = ~a + 1;
    for 

endmodule